`timescale 1ns / 1ps
`default_nettype none
//comment here
module update_wheel_tb();
  logic rst_in;

  logic clk_in;
  
  parameter POSITION_SIZE = 8;
  parameter VELOCITY_SIZE = 8;
  parameter NUM_VERTICES = 8;
  parameter NUM_OBSTACLES = 3;
  parameter NUM_NODES = 4;
  parameter NUM_SPRINGS = 6;
  parameter DT = 1;
  parameter ACCELERATION_SIZE = 8;
  parameter FORCE_SIZE = 8;
  parameter GRAVITY = -1;
  parameter TORQUE = 4;

  logic begin_update, result_out;
  logic [2:0] drive = 0;
  logic [$clog2(NUM_NODES)-1:0] springs [1:0][NUM_SPRINGS];
  logic signed [POSITION_SIZE-1:0] ideal [1:0][NUM_NODES];
  logic signed [POSITION_SIZE-1:0] obstacles [1:0][NUM_VERTICES][NUM_OBSTACLES];
  logic [$clog2(NUM_VERTICES):0] all_num_vertices [NUM_OBSTACLES];
  logic [POSITION_SIZE-1:0] axle [1:0];
  logic [$clog2(NUM_OBSTACLES)-1:0] num_obstacles;
  logic signed [POSITION_SIZE-1:0] nodes [1:0][NUM_NODES];
  logic signed [VELOCITY_SIZE-1:0] velocities [1:0][NUM_NODES];
  logic signed [FORCE_SIZE-1:0] axle_force [1:0];
  logic signed [VELOCITY_SIZE-1:0] axle_velocity [1:0];
  //logic signed [POSITION_SIZE-1:0] com [1:0];

  assign axle[0] = 5;
  assign axle[1] = 2;
  assign axle_velocity[0] = 0;
  assign axle_velocity[1] = 0;
  //obstacles must be oriented clockwise
  //obstacle 1
  assign obstacles[0][0][0] = -10; //point 1
  assign obstacles[1][0][0] = -10;        
  assign obstacles[0][1][0] = 10; //point 2
  assign obstacles[1][1][0] = -10;  
  assign obstacles[0][2][0] = 10;  //point 3
  assign obstacles[1][2][0] = 10;
  assign obstacles[0][3][0] = 15;  //point 4
  assign obstacles[1][3][0] = 10;
  assign obstacles[0][4][0] = 15;  //point 5
  assign obstacles[1][4][0] = -15;
  assign obstacles[0][5][0] = -15;  //point 6
  assign obstacles[1][5][0] = -15;
  assign obstacles[0][6][0] = -15;  //point 7
  assign obstacles[1][6][0] = 10;
  assign obstacles[0][7][0] = -10;  //point 8
  assign obstacles[1][7][0] = 10;

  assign all_num_vertices[0] = 8;
  assign num_obstacles = 1;

  assign nodes[0][0] = -3;
  assign nodes[1][0] = -2;
  assign nodes[0][1] = -2;
  assign nodes[1][1] = 2;
  assign nodes[0][2] = 2;
  assign nodes[1][2] = 2;
  assign nodes[0][3] = 3;
  assign nodes[1][3] = -2;

  assign ideal[0][0] = -3;
  assign ideal[1][0] = -2;
  assign ideal[0][1] = -2;
  assign ideal[1][1] = 2;
  assign ideal[0][2] = 2;
  assign ideal[1][2] = 2;
  assign ideal[0][3] = 3;
  assign ideal[1][3] = -2;

  assign springs[0][0] = 0;
  assign springs[1][0] = 1;
  assign springs[0][1] = 1;
  assign springs[1][1] = 2;
  assign springs[0][2] = 2;
  assign springs[1][2] = 3;
  assign springs[0][3] = 3;
  assign springs[1][3] = 0;
  assign springs[0][4] = 0;
  assign springs[1][4] = 2;
  assign springs[0][5] = 1;
  assign springs[1][5] = 3;

  assign velocities[0][0] = 0;
  assign velocities[1][0] = 0;
  assign velocities[0][1] = 0;
  assign velocities[1][1] = 0;
  assign velocities[0][2] = 0;
  assign velocities[1][2] = 0;
  assign velocities[0][3] = 0;
  assign velocities[1][3] = 0;

  // Instantiate the update_wheel module
  update_wheel #(
    .NUM_SPRINGS(NUM_SPRINGS),
    .NUM_NODES(NUM_NODES),
    .NUM_VERTICES(NUM_VERTICES),
    .NUM_OBSTACLES(NUM_OBSTACLES),
    .POSITION_SIZE(POSITION_SIZE),
    .VELOCITY_SIZE(VELOCITY_SIZE),
    .FORCE_SIZE(FORCE_SIZE),
    .TORQUE(TORQUE),
    .GRAVITY(GRAVITY),
    .DT(DT)
  ) wheel_updater (
    .clk_in(clk_in),
    .rst_in(rst_in),
    .begin_in(begin_update),
    .drive(drive),
    .ideal(ideal),
    .obstacles(obstacles),
    .all_num_vertices(all_num_vertices),
    .num_obstacles(num_obstacles),
    .nodes_in(nodes),
    .velocities_in(velocities),
    .springs(springs),
    .axle(axle),
    .axle_velocity(axle_velocity),
    .nodes_out(new_nodes),
    .velocities_out(new_velocities),
    .axle_force(axle_force),
    .result_out(result_out)
  );

  logic signed [POSITION_SIZE-1:0] new_nodes [1:0][NUM_NODES];
  logic signed [VELOCITY_SIZE-1:0] new_velocities [1:0][NUM_NODES];
  //logic signed [POSITION_SIZE-1:0] new_com [1:0];

  always begin
      #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
      clk_in = !clk_in;
  end
  always begin
    #10
    if (result_out == 1) begin
      begin_update <= 1;
      #10
      begin_update <= 0;
    end
        
  end
  //initial block...this is our test simulation
  initial begin
    $dumpfile("vsg.vcd"); //file to store value change dump (vcd)
    $dumpvars(1,update_wheel_tb,wheel_updater,wheel_updater.collider, wheel_updater.collider.collision_doer, wheel_updater.ideal_instance, wheel_updater.ideal_instance.springs_instance);

    $display("Starting Sim"); //print nice message at start
    clk_in = 1;
    rst_in = 0;
    #10;
    rst_in = 1;
    #10;
    rst_in = 0;
    begin_update = 1;
    #10
    begin_update = 0;

    #30000

    $display("Simulation finished");
    $finish;
  end
endmodule
`default_nettype wire